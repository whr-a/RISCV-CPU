`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/10/30 15:30:44
// Design Name: 
// Module Name: iFetch
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`ifndef IFETCH
`define IFETCH
`include "SetSize.v"
module iFetch(
    input wire clk,
    input wire rst,
    input wire rdy
     
    );
endmodule
`endif